library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity wfmlut is
	port (
		addr : in std_logic_vector (7 downto 0);
		sin  : out std_logic_vector (15 downto 0);
		cos  : out std_logic_vector (15 downto 0)
	);
end entity;

architecture arch of wfmlut is
begin

	process (addr)
	begin
		case addr is
			when "00000000" => sin <= "0000000000000000"; cos <= "0111111111111111";
			when "00000001" => sin <= "0000001100100100"; cos <= "0111111111110110";
			when "00000010" => sin <= "0000011001001000"; cos <= "0111111111011001";
			when "00000011" => sin <= "0000100101101011"; cos <= "0111111110100111";
			when "00000100" => sin <= "0000110010001100"; cos <= "0111111101100010";
			when "00000101" => sin <= "0000111110101011"; cos <= "0111111100001010";
			when "00000110" => sin <= "0001001011001000"; cos <= "0111111010011101";
			when "00000111" => sin <= "0001010111100010"; cos <= "0111111000011110";
			when "00001000" => sin <= "0001100011111001"; cos <= "0111110110001010";
			when "00001001" => sin <= "0001110000001100"; cos <= "0111110011100100";
			when "00001010" => sin <= "0001111100011010"; cos <= "0111110000101010";
			when "00001011" => sin <= "0010001000100100"; cos <= "0111101101011101";
			when "00001100" => sin <= "0010010100101000"; cos <= "0111101001111101";
			when "00001101" => sin <= "0010100000100111"; cos <= "0111100110001010";
			when "00001110" => sin <= "0010101100011111"; cos <= "0111100010000101";
			when "00001111" => sin <= "0010111000010001"; cos <= "0111011101101100";
			when "00010000" => sin <= "0011000011111100"; cos <= "0111011001000010";
			when "00010001" => sin <= "0011001111011111"; cos <= "0111010100000101";
			when "00010010" => sin <= "0011011010111010"; cos <= "0111001110110110";
			when "00010011" => sin <= "0011100110001101"; cos <= "0111001001010101";
			when "00010100" => sin <= "0011110001010111"; cos <= "0111000011100011";
			when "00010101" => sin <= "0011111100010111"; cos <= "0110111101011111";
			when "00010110" => sin <= "0100000111001110"; cos <= "0110110111001010";
			when "00010111" => sin <= "0100010001111011"; cos <= "0110110000100100";
			when "00011000" => sin <= "0100011100011101"; cos <= "0110101001101110";
			when "00011001" => sin <= "0100100110110100"; cos <= "0110100010100111";
			when "00011010" => sin <= "0100110001000000"; cos <= "0110011011010000";
			when "00011011" => sin <= "0100111011000000"; cos <= "0110010011101001";
			when "00011100" => sin <= "0101000100110100"; cos <= "0110001011110010";
			when "00011101" => sin <= "0101001110011011"; cos <= "0110000011101100";
			when "00011110" => sin <= "0101010111110110"; cos <= "0101111011010111";
			when "00011111" => sin <= "0101100001000011"; cos <= "0101110010110100";
			when "00100000" => sin <= "0101101010000010"; cos <= "0101101010000010";
			when "00100001" => sin <= "0101110010110100"; cos <= "0101100001000011";
			when "00100010" => sin <= "0101111011010111"; cos <= "0101010111110110";
			when "00100011" => sin <= "0110000011101100"; cos <= "0101001110011011";
			when "00100100" => sin <= "0110001011110010"; cos <= "0101000100110100";
			when "00100101" => sin <= "0110010011101001"; cos <= "0100111011000000";
			when "00100110" => sin <= "0110011011010000"; cos <= "0100110001000000";
			when "00100111" => sin <= "0110100010100111"; cos <= "0100100110110100";
			when "00101000" => sin <= "0110101001101110"; cos <= "0100011100011101";
			when "00101001" => sin <= "0110110000100100"; cos <= "0100010001111011";
			when "00101010" => sin <= "0110110111001010"; cos <= "0100000111001110";
			when "00101011" => sin <= "0110111101011111"; cos <= "0011111100010111";
			when "00101100" => sin <= "0111000011100011"; cos <= "0011110001010111";
			when "00101101" => sin <= "0111001001010101"; cos <= "0011100110001101";
			when "00101110" => sin <= "0111001110110110"; cos <= "0011011010111010";
			when "00101111" => sin <= "0111010100000101"; cos <= "0011001111011111";
			when "00110000" => sin <= "0111011001000010"; cos <= "0011000011111100";
			when "00110001" => sin <= "0111011101101100"; cos <= "0010111000010001";
			when "00110010" => sin <= "0111100010000101"; cos <= "0010101100011111";
			when "00110011" => sin <= "0111100110001010"; cos <= "0010100000100111";
			when "00110100" => sin <= "0111101001111101"; cos <= "0010010100101000";
			when "00110101" => sin <= "0111101101011101"; cos <= "0010001000100100";
			when "00110110" => sin <= "0111110000101010"; cos <= "0001111100011010";
			when "00110111" => sin <= "0111110011100100"; cos <= "0001110000001100";
			when "00111000" => sin <= "0111110110001010"; cos <= "0001100011111001";
			when "00111001" => sin <= "0111111000011110"; cos <= "0001010111100010";
			when "00111010" => sin <= "0111111010011101"; cos <= "0001001011001000";
			when "00111011" => sin <= "0111111100001010"; cos <= "0000111110101011";
			when "00111100" => sin <= "0111111101100010"; cos <= "0000110010001100";
			when "00111101" => sin <= "0111111110100111"; cos <= "0000100101101011";
			when "00111110" => sin <= "0111111111011001"; cos <= "0000011001001000";
			when "00111111" => sin <= "0111111111110110"; cos <= "0000001100100100";
			when "01000000" => sin <= "0111111111111111"; cos <= "0000000000000000";
			when "01000001" => sin <= "0111111111110110"; cos <= "1111110011011100";
			when "01000010" => sin <= "0111111111011001"; cos <= "1111100110111000";
			when "01000011" => sin <= "0111111110100111"; cos <= "1111011010010101";
			when "01000100" => sin <= "0111111101100010"; cos <= "1111001101110100";
			when "01000101" => sin <= "0111111100001010"; cos <= "1111000001010101";
			when "01000110" => sin <= "0111111010011101"; cos <= "1110110100111000";
			when "01000111" => sin <= "0111111000011110"; cos <= "1110101000011110";
			when "01001000" => sin <= "0111110110001010"; cos <= "1110011100000111";
			when "01001001" => sin <= "0111110011100100"; cos <= "1110001111110100";
			when "01001010" => sin <= "0111110000101010"; cos <= "1110000011100110";
			when "01001011" => sin <= "0111101101011101"; cos <= "1101110111011100";
			when "01001100" => sin <= "0111101001111101"; cos <= "1101101011011000";
			when "01001101" => sin <= "0111100110001010"; cos <= "1101011111011001";
			when "01001110" => sin <= "0111100010000101"; cos <= "1101010011100001";
			when "01001111" => sin <= "0111011101101100"; cos <= "1101000111101111";
			when "01010000" => sin <= "0111011001000010"; cos <= "1100111100000100";
			when "01010001" => sin <= "0111010100000101"; cos <= "1100110000100001";
			when "01010010" => sin <= "0111001110110110"; cos <= "1100100101000110";
			when "01010011" => sin <= "0111001001010101"; cos <= "1100011001110011";
			when "01010100" => sin <= "0111000011100011"; cos <= "1100001110101001";
			when "01010101" => sin <= "0110111101011111"; cos <= "1100000011101001";
			when "01010110" => sin <= "0110110111001010"; cos <= "1011111000110010";
			when "01010111" => sin <= "0110110000100100"; cos <= "1011101110000101";
			when "01011000" => sin <= "0110101001101110"; cos <= "1011100011100011";
			when "01011001" => sin <= "0110100010100111"; cos <= "1011011001001100";
			when "01011010" => sin <= "0110011011010000"; cos <= "1011001111000000";
			when "01011011" => sin <= "0110010011101001"; cos <= "1011000101000000";
			when "01011100" => sin <= "0110001011110010"; cos <= "1010111011001100";
			when "01011101" => sin <= "0110000011101100"; cos <= "1010110001100101";
			when "01011110" => sin <= "0101111011010111"; cos <= "1010101000001010";
			when "01011111" => sin <= "0101110010110100"; cos <= "1010011110111101";
			when "01100000" => sin <= "0101101010000010"; cos <= "1010010101111110";
			when "01100001" => sin <= "0101100001000011"; cos <= "1010001101001100";
			when "01100010" => sin <= "0101010111110110"; cos <= "1010000100101001";
			when "01100011" => sin <= "0101001110011011"; cos <= "1001111100010100";
			when "01100100" => sin <= "0101000100110100"; cos <= "1001110100001110";
			when "01100101" => sin <= "0100111011000000"; cos <= "1001101100010111";
			when "01100110" => sin <= "0100110001000000"; cos <= "1001100100110000";
			when "01100111" => sin <= "0100100110110100"; cos <= "1001011101011001";
			when "01101000" => sin <= "0100011100011101"; cos <= "1001010110010010";
			when "01101001" => sin <= "0100010001111011"; cos <= "1001001111011100";
			when "01101010" => sin <= "0100000111001110"; cos <= "1001001000110110";
			when "01101011" => sin <= "0011111100010111"; cos <= "1001000010100001";
			when "01101100" => sin <= "0011110001010111"; cos <= "1000111100011101";
			when "01101101" => sin <= "0011100110001101"; cos <= "1000110110101011";
			when "01101110" => sin <= "0011011010111010"; cos <= "1000110001001010";
			when "01101111" => sin <= "0011001111011111"; cos <= "1000101011111011";
			when "01110000" => sin <= "0011000011111100"; cos <= "1000100110111110";
			when "01110001" => sin <= "0010111000010001"; cos <= "1000100010010100";
			when "01110010" => sin <= "0010101100011111"; cos <= "1000011101111011";
			when "01110011" => sin <= "0010100000100111"; cos <= "1000011001110110";
			when "01110100" => sin <= "0010010100101000"; cos <= "1000010110000011";
			when "01110101" => sin <= "0010001000100100"; cos <= "1000010010100011";
			when "01110110" => sin <= "0001111100011010"; cos <= "1000001111010110";
			when "01110111" => sin <= "0001110000001100"; cos <= "1000001100011100";
			when "01111000" => sin <= "0001100011111001"; cos <= "1000001001110110";
			when "01111001" => sin <= "0001010111100010"; cos <= "1000000111100010";
			when "01111010" => sin <= "0001001011001000"; cos <= "1000000101100011";
			when "01111011" => sin <= "0000111110101011"; cos <= "1000000011110110";
			when "01111100" => sin <= "0000110010001100"; cos <= "1000000010011110";
			when "01111101" => sin <= "0000100101101011"; cos <= "1000000001011001";
			when "01111110" => sin <= "0000011001001000"; cos <= "1000000000100111";
			when "01111111" => sin <= "0000001100100100"; cos <= "1000000000001010";
			when "10000000" => sin <= "0000000000000000"; cos <= "1000000000000000";
			when "10000001" => sin <= "1111110011011100"; cos <= "1000000000001010";
			when "10000010" => sin <= "1111100110111000"; cos <= "1000000000100111";
			when "10000011" => sin <= "1111011010010101"; cos <= "1000000001011001";
			when "10000100" => sin <= "1111001101110100"; cos <= "1000000010011110";
			when "10000101" => sin <= "1111000001010101"; cos <= "1000000011110110";
			when "10000110" => sin <= "1110110100111000"; cos <= "1000000101100011";
			when "10000111" => sin <= "1110101000011110"; cos <= "1000000111100010";
			when "10001000" => sin <= "1110011100000111"; cos <= "1000001001110110";
			when "10001001" => sin <= "1110001111110100"; cos <= "1000001100011100";
			when "10001010" => sin <= "1110000011100110"; cos <= "1000001111010110";
			when "10001011" => sin <= "1101110111011100"; cos <= "1000010010100011";
			when "10001100" => sin <= "1101101011011000"; cos <= "1000010110000011";
			when "10001101" => sin <= "1101011111011001"; cos <= "1000011001110110";
			when "10001110" => sin <= "1101010011100001"; cos <= "1000011101111011";
			when "10001111" => sin <= "1101000111101111"; cos <= "1000100010010100";
			when "10010000" => sin <= "1100111100000100"; cos <= "1000100110111110";
			when "10010001" => sin <= "1100110000100001"; cos <= "1000101011111011";
			when "10010010" => sin <= "1100100101000110"; cos <= "1000110001001010";
			when "10010011" => sin <= "1100011001110011"; cos <= "1000110110101011";
			when "10010100" => sin <= "1100001110101001"; cos <= "1000111100011101";
			when "10010101" => sin <= "1100000011101001"; cos <= "1001000010100001";
			when "10010110" => sin <= "1011111000110010"; cos <= "1001001000110110";
			when "10010111" => sin <= "1011101110000101"; cos <= "1001001111011100";
			when "10011000" => sin <= "1011100011100011"; cos <= "1001010110010010";
			when "10011001" => sin <= "1011011001001100"; cos <= "1001011101011001";
			when "10011010" => sin <= "1011001111000000"; cos <= "1001100100110000";
			when "10011011" => sin <= "1011000101000000"; cos <= "1001101100010111";
			when "10011100" => sin <= "1010111011001100"; cos <= "1001110100001110";
			when "10011101" => sin <= "1010110001100101"; cos <= "1001111100010100";
			when "10011110" => sin <= "1010101000001010"; cos <= "1010000100101001";
			when "10011111" => sin <= "1010011110111101"; cos <= "1010001101001100";
			when "10100000" => sin <= "1010010101111110"; cos <= "1010010101111110";
			when "10100001" => sin <= "1010001101001100"; cos <= "1010011110111101";
			when "10100010" => sin <= "1010000100101001"; cos <= "1010101000001010";
			when "10100011" => sin <= "1001111100010100"; cos <= "1010110001100101";
			when "10100100" => sin <= "1001110100001110"; cos <= "1010111011001100";
			when "10100101" => sin <= "1001101100010111"; cos <= "1011000101000000";
			when "10100110" => sin <= "1001100100110000"; cos <= "1011001111000000";
			when "10100111" => sin <= "1001011101011001"; cos <= "1011011001001100";
			when "10101000" => sin <= "1001010110010010"; cos <= "1011100011100011";
			when "10101001" => sin <= "1001001111011100"; cos <= "1011101110000101";
			when "10101010" => sin <= "1001001000110110"; cos <= "1011111000110010";
			when "10101011" => sin <= "1001000010100001"; cos <= "1100000011101001";
			when "10101100" => sin <= "1000111100011101"; cos <= "1100001110101001";
			when "10101101" => sin <= "1000110110101011"; cos <= "1100011001110011";
			when "10101110" => sin <= "1000110001001010"; cos <= "1100100101000110";
			when "10101111" => sin <= "1000101011111011"; cos <= "1100110000100001";
			when "10110000" => sin <= "1000100110111110"; cos <= "1100111100000100";
			when "10110001" => sin <= "1000100010010100"; cos <= "1101000111101111";
			when "10110010" => sin <= "1000011101111011"; cos <= "1101010011100001";
			when "10110011" => sin <= "1000011001110110"; cos <= "1101011111011001";
			when "10110100" => sin <= "1000010110000011"; cos <= "1101101011011000";
			when "10110101" => sin <= "1000010010100011"; cos <= "1101110111011100";
			when "10110110" => sin <= "1000001111010110"; cos <= "1110000011100110";
			when "10110111" => sin <= "1000001100011100"; cos <= "1110001111110100";
			when "10111000" => sin <= "1000001001110110"; cos <= "1110011100000111";
			when "10111001" => sin <= "1000000111100010"; cos <= "1110101000011110";
			when "10111010" => sin <= "1000000101100011"; cos <= "1110110100111000";
			when "10111011" => sin <= "1000000011110110"; cos <= "1111000001010101";
			when "10111100" => sin <= "1000000010011110"; cos <= "1111001101110100";
			when "10111101" => sin <= "1000000001011001"; cos <= "1111011010010101";
			when "10111110" => sin <= "1000000000100111"; cos <= "1111100110111000";
			when "10111111" => sin <= "1000000000001010"; cos <= "1111110011011100";
			when "11000000" => sin <= "1000000000000000"; cos <= "0000000000000000";
			when "11000001" => sin <= "1000000000001010"; cos <= "0000001100100100";
			when "11000010" => sin <= "1000000000100111"; cos <= "0000011001001000";
			when "11000011" => sin <= "1000000001011001"; cos <= "0000100101101011";
			when "11000100" => sin <= "1000000010011110"; cos <= "0000110010001100";
			when "11000101" => sin <= "1000000011110110"; cos <= "0000111110101011";
			when "11000110" => sin <= "1000000101100011"; cos <= "0001001011001000";
			when "11000111" => sin <= "1000000111100010"; cos <= "0001010111100010";
			when "11001000" => sin <= "1000001001110110"; cos <= "0001100011111001";
			when "11001001" => sin <= "1000001100011100"; cos <= "0001110000001100";
			when "11001010" => sin <= "1000001111010110"; cos <= "0001111100011010";
			when "11001011" => sin <= "1000010010100011"; cos <= "0010001000100100";
			when "11001100" => sin <= "1000010110000011"; cos <= "0010010100101000";
			when "11001101" => sin <= "1000011001110110"; cos <= "0010100000100111";
			when "11001110" => sin <= "1000011101111011"; cos <= "0010101100011111";
			when "11001111" => sin <= "1000100010010100"; cos <= "0010111000010001";
			when "11010000" => sin <= "1000100110111110"; cos <= "0011000011111100";
			when "11010001" => sin <= "1000101011111011"; cos <= "0011001111011111";
			when "11010010" => sin <= "1000110001001010"; cos <= "0011011010111010";
			when "11010011" => sin <= "1000110110101011"; cos <= "0011100110001101";
			when "11010100" => sin <= "1000111100011101"; cos <= "0011110001010111";
			when "11010101" => sin <= "1001000010100001"; cos <= "0011111100010111";
			when "11010110" => sin <= "1001001000110110"; cos <= "0100000111001110";
			when "11010111" => sin <= "1001001111011100"; cos <= "0100010001111011";
			when "11011000" => sin <= "1001010110010010"; cos <= "0100011100011101";
			when "11011001" => sin <= "1001011101011001"; cos <= "0100100110110100";
			when "11011010" => sin <= "1001100100110000"; cos <= "0100110001000000";
			when "11011011" => sin <= "1001101100010111"; cos <= "0100111011000000";
			when "11011100" => sin <= "1001110100001110"; cos <= "0101000100110100";
			when "11011101" => sin <= "1001111100010100"; cos <= "0101001110011011";
			when "11011110" => sin <= "1010000100101001"; cos <= "0101010111110110";
			when "11011111" => sin <= "1010001101001100"; cos <= "0101100001000011";
			when "11100000" => sin <= "1010010101111110"; cos <= "0101101010000010";
			when "11100001" => sin <= "1010011110111101"; cos <= "0101110010110100";
			when "11100010" => sin <= "1010101000001010"; cos <= "0101111011010111";
			when "11100011" => sin <= "1010110001100101"; cos <= "0110000011101100";
			when "11100100" => sin <= "1010111011001100"; cos <= "0110001011110010";
			when "11100101" => sin <= "1011000101000000"; cos <= "0110010011101001";
			when "11100110" => sin <= "1011001111000000"; cos <= "0110011011010000";
			when "11100111" => sin <= "1011011001001100"; cos <= "0110100010100111";
			when "11101000" => sin <= "1011100011100011"; cos <= "0110101001101110";
			when "11101001" => sin <= "1011101110000101"; cos <= "0110110000100100";
			when "11101010" => sin <= "1011111000110010"; cos <= "0110110111001010";
			when "11101011" => sin <= "1100000011101001"; cos <= "0110111101011111";
			when "11101100" => sin <= "1100001110101001"; cos <= "0111000011100011";
			when "11101101" => sin <= "1100011001110011"; cos <= "0111001001010101";
			when "11101110" => sin <= "1100100101000110"; cos <= "0111001110110110";
			when "11101111" => sin <= "1100110000100001"; cos <= "0111010100000101";
			when "11110000" => sin <= "1100111100000100"; cos <= "0111011001000010";
			when "11110001" => sin <= "1101000111101111"; cos <= "0111011101101100";
			when "11110010" => sin <= "1101010011100001"; cos <= "0111100010000101";
			when "11110011" => sin <= "1101011111011001"; cos <= "0111100110001010";
			when "11110100" => sin <= "1101101011011000"; cos <= "0111101001111101";
			when "11110101" => sin <= "1101110111011100"; cos <= "0111101101011101";
			when "11110110" => sin <= "1110000011100110"; cos <= "0111110000101010";
			when "11110111" => sin <= "1110001111110100"; cos <= "0111110011100100";
			when "11111000" => sin <= "1110011100000111"; cos <= "0111110110001010";
			when "11111001" => sin <= "1110101000011110"; cos <= "0111111000011110";
			when "11111010" => sin <= "1110110100111000"; cos <= "0111111010011101";
			when "11111011" => sin <= "1111000001010101"; cos <= "0111111100001010";
			when "11111100" => sin <= "1111001101110100"; cos <= "0111111101100010";
			when "11111101" => sin <= "1111011010010101"; cos <= "0111111110100111";
			when "11111110" => sin <= "1111100110111000"; cos <= "0111111111011001";
			when "11111111" => sin <= "1111110011011100"; cos <= "0111111111110110";
			when others => sin <= (others => '0'); cos <= (others => '0');
		end case;
	end process;

end architecture;
